ENTITY and_3 IS
	PORT (a,b,c: IN bit; output: OUT bit);	
END and_3;

ARCHITECTURE data_flow OF and_3 IS
BEGIN
	output <= a and b AND c;
END data_flow;
		