ENTITY or_5 IS
	PORT(a,b,c,d,e: IN bit; output: OUT bit);
END or_5;

ARCHITECTURE data_flow OF or_5 IS
BEGIN
	output <= a OR b OR c OR d OR e;
END data_flow;